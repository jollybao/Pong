----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:25:49 03/03/2016 
-- Design Name: 
-- Module Name:    font_rom - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity font_rom is
	port(
		addr: in std_logic_vector(10 downto 0);
		dataOut: out std_logic_vector(7 downto 0)
	);
end font_rom;

architecture Behavioral of font_rom is
   
	signal data: STD_LOGIC_VECTOR(7 downto 0);
	type rom_type is array (0 to 2047) of std_logic_vector(0 to 7);

	-- ROM definition
	constant ROM: rom_type := (   -- 2^11-by-8
		-- NUL: code x00
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- SOH: code x01
		"00000000", -- 0
		"00000000", -- 1
		"01111110", -- 2  ******
		"10000001", -- 3 *      *
		"10100101", -- 4 * *  * *
		"10000001", -- 5 *      *
		"10000001", -- 6 *      *
		"10111101", -- 7 * **** *
		"10011001", -- 8 *  **  *
		"10000001", -- 9 *      *
		"10000001", -- a *      *
		"01111110", -- b  ******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- STX: code x02
		"00000000", -- 0
		"00000000", -- 1
		"01111110", -- 2  ******
		"11111111", -- 3 ********
		"11011011", -- 4 ** ** **
		"11111111", -- 5 ********
		"11111111", -- 6 ********
		"11000011", -- 7 **    **
		"11100111", -- 8 ***  ***
		"11111111", -- 9 ********
		"11111111", -- a ********
		"01111110", -- b  ******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- ETX: code x03
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"01101100", -- 4  ** **
		"11111110", -- 5 *******
		"11111110", -- 6 *******
		"11111110", -- 7 *******
		"11111110", -- 8 *******
		"01111100", -- 9  *****
		"00111000", -- a   ***
		"00010000", -- b    *
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- EOT: code x04
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00010000", -- 4    *
		"00111000", -- 5   ***
		"01111100", -- 6  *****
		"11111110", -- 7 *******
		"01111100", -- 8  *****
		"00111000", -- 9   ***
		"00010000", -- a    *
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- ENQ: code x05
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00011000", -- 3    **
		"00111100", -- 4   ****
		"00111100", -- 5   ****
		"11100111", -- 6 ***  ***
		"11100111", -- 7 ***  ***
		"11100111", -- 8 ***  ***
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- ACK: code x06
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00011000", -- 3    **
		"00111100", -- 4   ****
		"01111110", -- 5  ******
		"11111111", -- 6 ********
		"11111111", -- 7 ********
		"01111110", -- 8  ******
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- BEL: code x07
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00011000", -- 6    **
		"00111100", -- 7   ****
		"00111100", -- 8   ****
		"00011000", -- 9    **
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- BS: code x08
		"11111111", -- 0 ********
		"11111111", -- 1 ********
		"11111111", -- 2 ********
		"11111111", -- 3 ********
		"11111111", -- 4 ********
		"11111111", -- 5 ********
		"11100111", -- 6 ***  ***
		"11000011", -- 7 **    **
		"11000011", -- 8 **    **
		"11100111", -- 9 ***  ***
		"11111111", -- a ********
		"11111111", -- b ********
		"11111111", -- c ********
		"11111111", -- d ********
		"11111111", -- e ********
		"11111111", -- f ********
		-- HT: code x09
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00111100", -- 5   ****
		"01100110", -- 6  **  **
		"01000010", -- 7  *    *
		"01000010", -- 8  *    *
		"01100110", -- 9  **  **
		"00111100", -- a   ****
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- LF: code x0a
		"11111111", -- 0 ********
		"11111111", -- 1 ********
		"11111111", -- 2 ********
		"11111111", -- 3 ********
		"11111111", -- 4 ********
		"11000011", -- 5 **    **
		"10011001", -- 6 *  **  *
		"10111101", -- 7 * **** *
		"10111101", -- 8 * **** *
		"10011001", -- 9 *  **  *
		"11000011", -- a **    **
		"11111111", -- b ********
		"11111111", -- c ********
		"11111111", -- d ********
		"11111111", -- e ********
		"11111111", -- f ********
		-- code x0b
		"00000000", -- 0
		"00000000", -- 1
		"00011110", -- 2    ****
		"00001110", -- 3     ***
		"00011010", -- 4    ** *
		"00110010", -- 5   **  *
		"01111000", -- 6  ****
		"11001100", -- 7 **  **
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01111000", -- b  ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x0c
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01100110", -- 6  **  **
		"00111100", -- 7   ****
		"00011000", -- 8    **
		"01111110", -- 9  ******
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x0d
		"00000000", -- 0
		"00000000", -- 1
		"00111111", -- 2   ******
		"00110011", -- 3   **  **
		"00111111", -- 4   ******
		"00110000", -- 5   **
		"00110000", -- 6   **
		"00110000", -- 7   **
		"00110000", -- 8   **
		"01110000", -- 9  ***
		"11110000", -- a ****
		"11100000", -- b ***
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x0e
		"00000000", -- 0
		"00000000", -- 1
		"01111111", -- 2  *******
		"01100011", -- 3  **   **
		"01111111", -- 4  *******
		"01100011", -- 5  **   **
		"01100011", -- 6  **   **
		"01100011", -- 7  **   **
		"01100011", -- 8  **   **
		"01100111", -- 9  **  ***
		"11100111", -- a ***  ***
		"11100110", -- b ***  **
		"11000000", -- c **
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x0f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00011000", -- 3    **
		"00011000", -- 4    **
		"11011011", -- 5 ** ** **
		"00111100", -- 6   ****
		"11100111", -- 7 ***  ***
		"00111100", -- 8   ****
		"11011011", -- 9 ** ** **
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x10
		"00000000", -- 0
		"10000000", -- 1 *
		"11000000", -- 2 **
		"11100000", -- 3 ***
		"11110000", -- 4 ****
		"11111000", -- 5 *****
		"11111110", -- 6 *******
		"11111000", -- 7 *****
		"11110000", -- 8 ****
		"11100000", -- 9 ***
		"11000000", -- a **
		"10000000", -- b *
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x11
		"00000000", -- 0
		"00000010", -- 1       *
		"00000110", -- 2      **
		"00001110", -- 3     ***
		"00011110", -- 4    ****
		"00111110", -- 5   *****
		"11111110", -- 6 *******
		"00111110", -- 7   *****
		"00011110", -- 8    ****
		"00001110", -- 9     ***
		"00000110", -- a      **
		"00000010", -- b       *
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x12
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00111100", -- 3   ****
		"01111110", -- 4  ******
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"01111110", -- 8  ******
		"00111100", -- 9   ****
		"00011000", -- a    **
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x13
		"00000000", -- 0
		"00000000", -- 1
		"01100110", -- 2  **  **
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01100110", -- 6  **  **
		"01100110", -- 7  **  **
		"01100110", -- 8  **  **
		"00000000", -- 9
		"01100110", -- a  **  **
		"01100110", -- b  **  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x14
		"00000000", -- 0
		"00000000", -- 1
		"01111111", -- 2  *******
		"11011011", -- 3 ** ** **
		"11011011", -- 4 ** ** **
		"11011011", -- 5 ** ** **
		"01111011", -- 6  **** **
		"00011011", -- 7    ** **
		"00011011", -- 8    ** **
		"00011011", -- 9    ** **
		"00011011", -- a    ** **
		"00011011", -- b    ** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x15
		"00000000", -- 0
		"01111100", -- 1  *****
		"11000110", -- 2 **   **
		"01100000", -- 3  **
		"00111000", -- 4   ***
		"01101100", -- 5  ** **
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"01101100", -- 8  ** **
		"00111000", -- 9   ***
		"00001100", -- a     **
		"11000110", -- b **   **
		"01111100", -- c  *****
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x16
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"11111110", -- 8 *******
		"11111110", -- 9 *******
		"11111110", -- a *******
		"11111110", -- b *******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x17
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00111100", -- 3   ****
		"01111110", -- 4  ******
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"01111110", -- 8  ******
		"00111100", -- 9   ****
		"00011000", -- a    **
		"01111110", -- b  ******
		"00110000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x18
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00111100", -- 3   ****
		"01111110", -- 4  ******
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x19
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"01111110", -- 9  ******
		"00111100", -- a   ****
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x1a
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00011000", -- 5    **
		"00001100", -- 6     **
		"11111110", -- 7 *******
		"00001100", -- 8     **
		"00011000", -- 9    **
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x1b
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00110000", -- 5   **
		"01100000", -- 6  **
		"11111110", -- 7 *******
		"01100000", -- 8  **
		"00110000", -- 9   **
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x1c
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"11000000", -- 6 **
		"11000000", -- 7 **
		"11000000", -- 8 **
		"11111110", -- 9 *******
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x1d
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00100100", -- 5   *  *
		"01100110", -- 6  **  **
		"11111111", -- 7 ********
		"01100110", -- 8  **  **
		"00100100", -- 9   *  *
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x1e
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00010000", -- 4    *
		"00111000", -- 5   ***
		"00111000", -- 6   ***
		"01111100", -- 7  *****
		"01111100", -- 8  *****
		"11111110", -- 9 *******
		"11111110", -- a *******
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x1f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"11111110", -- 4 *******
		"11111110", -- 5 *******
		"01111100", -- 6  *****
		"01111100", -- 7  *****
		"00111000", -- 8   ***
		"00111000", -- 9   ***
		"00010000", -- a    *
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x20
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x21
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00111100", -- 3   ****
		"00111100", -- 4   ****
		"00111100", -- 5   ****
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00000000", -- 9
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x22
		"00000000", -- 0
		"01100110", -- 1  **  **
		"01100110", -- 2  **  **
		"01100110", -- 3  **  **
		"00100100", -- 4   *  *
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x23
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"01101100", -- 3  ** **
		"01101100", -- 4  ** **
		"11111110", -- 5 *******
		"01101100", -- 6  ** **
		"01101100", -- 7  ** **
		"01101100", -- 8  ** **
		"11111110", -- 9 *******
		"01101100", -- a  ** **
		"01101100", -- b  ** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x24
		"00011000", -- 0     **
		"00011000", -- 1     **
		"01111100", -- 2   *****
		"11000110", -- 3  **   **
		"11000010", -- 4  **    *
		"11000000", -- 5  **
		"01111100", -- 6   *****
		"00000110", -- 7       **
		"00000110", -- 8       **
		"10000110", -- 9  *    **
		"11000110", -- a  **   **
		"01111100", -- b   *****
		"00011000", -- c     **
		"00011000", -- d     **
		"00000000", -- e
		"00000000", -- f
		-- code x25
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"11000010", -- 4 **    *
		"11000110", -- 5 **   **
		"00001100", -- 6     **
		"00011000", -- 7    **
		"00110000", -- 8   **
		"01100000", -- 9  **
		"11000110", -- a **   **
		"10000110", -- b *    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x26
		"00000000", -- 0
		"00000000", -- 1
		"00111000", -- 2   ***
		"01101100", -- 3  ** **
		"01101100", -- 4  ** **
		"00111000", -- 5   ***
		"01110110", -- 6  *** **
		"11011100", -- 7 ** ***
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01110110", -- b  *** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x27
		"00000000", -- 0
		"00110000", -- 1   **
		"00110000", -- 2   **
		"00110000", -- 3   **
		"01100000", -- 4  **
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x28
		"00000000", -- 0
		"00000000", -- 1
		"00001100", -- 2     **
		"00011000", -- 3    **
		"00110000", -- 4   **
		"00110000", -- 5   **
		"00110000", -- 6   **
		"00110000", -- 7   **
		"00110000", -- 8   **
		"00110000", -- 9   **
		"00011000", -- a    **
		"00001100", -- b     **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x29
		"00000000", -- 0
		"00000000", -- 1
		"00110000", -- 2   **
		"00011000", -- 3    **
		"00001100", -- 4     **
		"00001100", -- 5     **
		"00001100", -- 6     **
		"00001100", -- 7     **
		"00001100", -- 8     **
		"00001100", -- 9     **
		"00011000", -- a    **
		"00110000", -- b   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x2a
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01100110", -- 5  **  **
		"00111100", -- 6   ****
		"11111111", -- 7 ********
		"00111100", -- 8   ****
		"01100110", -- 9  **  **
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x2b
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00011000", -- 5    **
		"00011000", -- 6    **
		"01111110", -- 7  ******
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x2c
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00011000", -- 9    **
		"00011000", -- a    **
		"00011000", -- b    **
		"00110000", -- c   **
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x2d
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"01111110", -- 7  ******
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x2e
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x2f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000010", -- 4       *
		"00000110", -- 5      **
		"00001100", -- 6     **
		"00011000", -- 7    **
		"00110000", -- 8   **
		"01100000", -- 9  **
		"11000000", -- a **
		"10000000", -- b *
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- 0: code x30
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11001110", -- 5 **  ***
		"11011110", -- 6 ** ****
		"11110110", -- 7 **** **
		"11100110", -- 8 ***  **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- 1: code x31
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2
		"00111000", -- 3
		"01111000", -- 4    **
		"00011000", -- 5   ***
		"00011000", -- 6  ****
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"01111110", -- b    **
		"00000000", -- c    **
		"00000000", -- d  ******
		"00000000", -- e
		"00000000", -- f
		-- 2: code x32
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"00000110", -- 4      **
		"00001100", -- 5     **
		"00011000", -- 6    **
		"00110000", -- 7   **
		"01100000", -- 8  **
		"11000000", -- 9 **
		"11000110", -- a **   **
		"11111110", -- b *******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- 3: code x33
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"00000110", -- 4      **
		"00000110", -- 5      **
		"00111100", -- 6   ****
		"00000110", -- 7      **
		"00000110", -- 8      **
		"00000110", -- 9      **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- 4: code x34
		"00000000", -- 0
		"00000000", -- 1
		"00001100", -- 2     **
		"00011100", -- 3    ***
		"00111100", -- 4   ****
		"01101100", -- 5  ** **
		"11001100", -- 6 **  **
		"11111110", -- 7 *******
		"00001100", -- 8     **
		"00001100", -- 9     **
		"00001100", -- a     **
		"00011110", -- b    ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x35
		"00000000", -- 0
		"00000000", -- 1
		"11111110", -- 2 *******
		"11000000", -- 3 **
		"11000000", -- 4 **
		"11000000", -- 5 **
		"11111100", -- 6 ******
		"00000110", -- 7      **
		"00000110", -- 8      **
		"00000110", -- 9      **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x36
		"00000000", -- 0
		"00000000", -- 1
		"00111000", -- 2   ***
		"01100000", -- 3  **
		"11000000", -- 4 **
		"11000000", -- 5 **
		"11111100", -- 6 ******
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x37
		"00000000", -- 0
		"00000000", -- 1
		"11111110", -- 2 *******
		"11000110", -- 3 **   **
		"00000110", -- 4      **
		"00000110", -- 5      **
		"00001100", -- 6     **
		"00011000", -- 7    **
		"00110000", -- 8   **
		"00110000", -- 9   **
		"00110000", -- a   **
		"00110000", -- b   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x38
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"01111100", -- 6  *****
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x39
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"01111110", -- 6  ******
		"00000110", -- 7      **
		"00000110", -- 8      **
		"00000110", -- 9      **
		"00001100", -- a     **
		"01111000", -- b  ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x3a
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00011000", -- 9    **
		"00011000", -- a    **
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x3b
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00011000", -- 9    **
		"00011000", -- a    **
		"00110000", -- b   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x3c
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000110", -- 3      **
		"00001100", -- 4     **
		"00011000", -- 5    **
		"00110000", -- 6   **
		"01100000", -- 7  **
		"00110000", -- 8   **
		"00011000", -- 9    **
		"00001100", -- a     **
		"00000110", -- b      **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x3d
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01111110", -- 5  ******
		"00000000", -- 6
		"00000000", -- 7
		"01111110", -- 8  ******
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x3e
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"01100000", -- 3  **
		"00110000", -- 4   **
		"00011000", -- 5    **
		"00001100", -- 6     **
		"00000110", -- 7      **
		"00001100", -- 8     **
		"00011000", -- 9    **
		"00110000", -- a   **
		"01100000", -- b  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x3f
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"00001100", -- 5     **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00000000", -- 9
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x40
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11011110", -- 6 ** ****
		"11011110", -- 7 ** ****
		"11011110", -- 8 ** ****
		"11011100", -- 9 ** ***
		"11000000", -- a **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- A: code x41
		"00000000", -- 0
		"00000000", -- 1
		"00010000", -- 2    *
		"00111000", -- 3   ***
		"01101100", -- 4  ** **
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"11111110", -- 7 *******
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"11000110", -- b **   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- B: code x42
		"00000000", -- 0
		"00000000", -- 1
		"11111100", -- 2 ******
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01111100", -- 6  *****
		"01100110", -- 7  **  **
		"01100110", -- 8  **  **
		"01100110", -- 9  **  **
		"01100110", -- a  **  **
		"11111100", -- b ******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- C: code x43
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"01100110", -- 3  **  **
		"11000010", -- 4 **    *
		"11000000", -- 5 **
		"11000000", -- 6 **
		"11000000", -- 7 **
		"11000000", -- 8 **
		"11000010", -- 9 **    *
		"01100110", -- a  **  **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- D: code x44
		"00000000", -- 0
		"00000000", -- 1
		"11111000", -- 2 *****
		"01101100", -- 3  ** **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01100110", -- 6  **  **
		"01100110", -- 7  **  **
		"01100110", -- 8  **  **
		"01100110", -- 9  **  **
		"01101100", -- a  ** **
		"11111000", -- b *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x45
		"00000000", -- 0
		"00000000", -- 1
		"11111110", -- 2 *******
		"01100110", -- 3  **  **
		"01100010", -- 4  **   *
		"01101000", -- 5  ** *
		"01111000", -- 6  ****
		"01101000", -- 7  ** *
		"01100000", -- 8  **
		"01100010", -- 9  **   *
		"01100110", -- a  **  **
		"11111110", -- b *******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x46
		"00000000", -- 0
		"00000000", -- 1
		"11111110", -- 2 *******
		"01100110", -- 3  **  **
		"01100010", -- 4  **   *
		"01101000", -- 5  ** *
		"01111000", -- 6  ****
		"01101000", -- 7  ** *
		"01100000", -- 8  **
		"01100000", -- 9  **
		"01100000", -- a  **
		"11110000", -- b ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x47
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"01100110", -- 3  **  **
		"11000010", -- 4 **    *
		"11000000", -- 5 **
		"11000000", -- 6 **
		"11011110", -- 7 ** ****
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"01100110", -- a  **  **
		"00111010", -- b   *** *
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- H: code x48
		"00000000", -- 0
		"00000000", -- 1
		"11000110", -- 2 **   **
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11111110", -- 6 *******
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"11000110", -- b **   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- I: code x49
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- J: code x4a
		"00000000", -- 0
		"00000000", -- 1
		"00011110", -- 2    ****
		"00001100", -- 3     **
		"00001100", -- 4     **
		"00001100", -- 5     **
		"00001100", -- 6     **
		"00001100", -- 7     **
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01111000", -- b  ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- K: code x4b
		"00000000", -- 0
		"00000000", -- 1
		"11100110", -- 2 ***  **
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01101100", -- 5  ** **
		"01111000", -- 6  ****
		"01111000", -- 7  ****
		"01101100", -- 8  ** **
		"01100110", -- 9  **  **
		"01100110", -- a  **  **
		"11100110", -- b ***  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- L: code x4c
		"00000000", -- 0
		"00000000", -- 1
		"11110000", -- 2 ****
		"01100000", -- 3  **
		"01100000", -- 4  **
		"01100000", -- 5  **
		"01100000", -- 6  **
		"01100000", -- 7  **
		"01100000", -- 8  **
		"01100010", -- 9  **   *
		"01100110", -- a  **  **
		"11111110", -- b *******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- M: code x4d
		"00000000", -- 0
		"00000000", -- 1
		"11000011", -- 2 **    **
		"11100111", -- 3 ***  ***
		"11111111", -- 4 ********
		"11111111", -- 5 ********
		"11011011", -- 6 ** ** **
		"11000011", -- 7 **    **
		"11000011", -- 8 **    **
		"11000011", -- 9 **    **
		"11000011", -- a **    **
		"11000011", -- b **    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- N: code x4e
		"00000000", -- 0
		"00000000", -- 1
		"11000110", -- 2 **   **
		"11100110", -- 3 ***  **
		"11110110", -- 4 **** **
		"11111110", -- 5 *******
		"11011110", -- 6 ** ****
		"11001110", -- 7 **  ***
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"11000110", -- b **   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- O: code x4f
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- P: code x50
		"00000000", -- 0
		"00000000", -- 1
		"11111100", -- 2 ******
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01111100", -- 6  *****
		"01100000", -- 7  **
		"01100000", -- 8  **
		"01100000", -- 9  **
		"01100000", -- a  **
		"11110000", -- b ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- Q: code x510
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11010110", -- 9 ** * **
		"11011110", -- a ** ****
		"01111100", -- b  *****
		"00001100", -- c     **
		"00001110", -- d     ***
		"00000000", -- e
		"00000000", -- f
		-- code x52
		"00000000", -- 0
		"00000000", -- 1
		"11111100", -- 2 ******
		"01100110", -- 3  **  **
		"01100110", -- 4  **  **
		"01100110", -- 5  **  **
		"01111100", -- 6  *****
		"01101100", -- 7  ** **
		"01100110", -- 8  **  **
		"01100110", -- 9  **  **
		"01100110", -- a  **  **
		"11100110", -- b ***  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x53
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"01100000", -- 5  **
		"00111000", -- 6   ***
		"00001100", -- 7     **
		"00000110", -- 8      **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x54
		"00000000", -- 0
		"00000000", -- 1
		"11111111", -- 2 ********
		"11011011", -- 3 ** ** **
		"10011001", -- 4 *  **  *
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x55
		"00000000", -- 0
		"00000000", -- 1
		"11000110", -- 2 **   **
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x56
		"00000000", -- 0
		"00000000", -- 1
		"11000011", -- 2 **    **
		"11000011", -- 3 **    **
		"11000011", -- 4 **    **
		"11000011", -- 5 **    **
		"11000011", -- 6 **    **
		"11000011", -- 7 **    **
		"11000011", -- 8 **    **
		"01100110", -- 9  **  **
		"00111100", -- a   ****
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x57
		"00000000", -- 0
		"00000000", -- 1
		"11000011", -- 2 **    **
		"11000011", -- 3 **    **
		"11000011", -- 4 **    **
		"11000011", -- 5 **    **
		"11000011", -- 6 **    **
		"11011011", -- 7 ** ** **
		"11011011", -- 8 ** ** **
		"11111111", -- 9 ********
		"01100110", -- a  **  **
		"01100110", -- b  **  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f

		-- code x58
		"00000000", -- 0
		"00000000", -- 1
		"11000011", -- 2 **    **
		"11000011", -- 3 **    **
		"01100110", -- 4  **  **
		"00111100", -- 5   ****
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00111100", -- 8   ****
		"01100110", -- 9  **  **
		"11000011", -- a **    **
		"11000011", -- b **    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x59
		"00000000", -- 0
		"00000000", -- 1
		"11000011", -- 2 **    **
		"11000011", -- 3 **    **
		"11000011", -- 4 **    **
		"01100110", -- 5  **  **
		"00111100", -- 6   ****
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x5a
		"00000000", -- 0
		"00000000", -- 1
		"11111111", -- 2 ********
		"11000011", -- 3 **    **
		"10000110", -- 4 *    **
		"00001100", -- 5     **
		"00011000", -- 6    **
		"00110000", -- 7   **
		"01100000", -- 8  **
		"11000001", -- 9 **     *
		"11000011", -- a **    **
		"11111111", -- b ********
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x5b
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"00110000", -- 3   **
		"00110000", -- 4   **
		"00110000", -- 5   **
		"00110000", -- 6   **
		"00110000", -- 7   **
		"00110000", -- 8   **
		"00110000", -- 9   **
		"00110000", -- a   **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x5c
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"10000000", -- 3 *
		"11000000", -- 4 **
		"11100000", -- 5 ***
		"01110000", -- 6  ***
		"00111000", -- 7   ***
		"00011100", -- 8    ***
		"00001110", -- 9     ***
		"00000110", -- a      **
		"00000010", -- b       *
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x5d
		"00000000", -- 0
		"00000000", -- 1
		"00111100", -- 2   ****
		"00001100", -- 3     **
		"00001100", -- 4     **
		"00001100", -- 5     **
		"00001100", -- 6     **
		"00001100", -- 7     **
		"00001100", -- 8     **
		"00001100", -- 9     **
		"00001100", -- a     **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x5e
		"00010000", -- 0    *
		"00111000", -- 1   ***
		"01101100", -- 2  ** **
		"11000110", -- 3 **   **
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x5f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"11111111", -- d ********
		"00000000", -- e
		"00000000", -- f
		-- code x60
		"00110000", -- 0   **
		"00110000", -- 1   **
		"00011000", -- 2    **
		"00000000", -- 3
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- a: code x61
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01111000", -- 5  ****
		"00001100", -- 6     **
		"01111100", -- 7  *****
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01110110", -- b  *** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- b: code x62
		"00000000", -- 0
		"00000000", -- 1
		"11100000", -- 2  ***
		"01100000", -- 3   **
		"01100000", -- 4   **
		"01111000", -- 5   ****
		"01101100", -- 6   ** **
		"01100110", -- 7   **  **
		"01100110", -- 8   **  **
		"01100110", -- 9   **  **
		"01100110", -- a   **  **
		"01111100", -- b   *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- c: code x63
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01111100", -- 5  *****
		"11000110", -- 6 **   **
		"11000000", -- 7 **
		"11000000", -- 8 **
		"11000000", -- 9 **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- d: code x64
		"00000000", -- 0
		"00000000", -- 1
		"00011100", -- 2    ***
		"00001100", -- 3     **
		"00001100", -- 4     **
		"00111100", -- 5   ****
		"01101100", -- 6  ** **
		"11001100", -- 7 **  **
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01110110", -- b  *** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- e: code x65
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01111100", -- 5  *****
		"11000110", -- 6 **   **
		"11111110", -- 7 *******
		"11000000", -- 8 **
		"11000000", -- 9 **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- f: code x66
		"00000000", -- 0
		"00000000", -- 1
		"00111000", -- 2   ***
		"01101100", -- 3  ** **
		"01100100", -- 4  **  *
		"01100000", -- 5  **
		"11110000", -- 6 ****
		"01100000", -- 7  **
		"01100000", -- 8  **
		"01100000", -- 9  **
		"01100000", -- a  **
		"11110000", -- b ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- g: code x67
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01110110", -- 5  *** **
		"11001100", -- 6 **  **
		"11001100", -- 7 **  **
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01111100", -- b  *****
		"00001100", -- c     **
		"11001100", -- d **  **
		"01111000", -- e  ****
		"00000000", -- f
		-- h: code x68
		"00000000", -- 0
		"00000000", -- 1
		"11100000", -- 2 ***
		"01100000", -- 3  **
		"01100000", -- 4  **
		"01101100", -- 5  ** **
		"01110110", -- 6  *** **
		"01100110", -- 7  **  **
		"01100110", -- 8  **  **
		"01100110", -- 9  **  **
		"01100110", -- a  **  **
		"11100110", -- b ***  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- i: code x69
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00011000", -- 3    **
		"00000000", -- 4
		"00111000", -- 5   ***
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- j: code x6a
		"00000000", -- 0
		"00000000", -- 1
		"00000110", -- 2      **
		"00000110", -- 3      **
		"00000000", -- 4
		"00001110", -- 5     ***
		"00000110", -- 6      **
		"00000110", -- 7      **
		"00000110", -- 8      **
		"00000110", -- 9      **
		"00000110", -- a      **
		"00000110", -- b      **
		"01100110", -- c  **  **
		"01100110", -- d  **  **
		"00111100", -- e   ****
		"00000000", -- f
		-- k: code x6b
		"00000000", -- 0
		"00000000", -- 1
		"11100000", -- 2 ***
		"01100000", -- 3  **
		"01100000", -- 4  **
		"01100110", -- 5  **  **
		"01101100", -- 6  ** **
		"01111000", -- 7  ****
		"01111000", -- 8  ****
		"01101100", -- 9  ** **
		"01100110", -- a  **  **
		"11100110", -- b ***  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- l: code x6c
		"00000000", -- 0
		"00000000", -- 1
		"00111000", -- 2   ***
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00011000", -- 6    **
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00111100", -- b   ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- m: code x6d
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11100110", -- 5 ***  **
		"11111111", -- 6 ********
		"11011011", -- 7 ** ** **
		"11011011", -- 8 ** ** **
		"11011011", -- 9 ** ** **
		"11011011", -- a ** ** **
		"11011011", -- b ** ** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- n: code x6e
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11011100", -- 5 ** ***
		"01100110", -- 6  **  **
		"01100110", -- 7  **  **
		"01100110", -- 8  **  **
		"01100110", -- 9  **  **
		"01100110", -- a  **  **
		"01100110", -- b  **  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- o: code x6f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01111100", -- 5  *****
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x70
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11011100", -- 5 ** ***
		"01100110", -- 6  **  **
		"01100110", -- 7  **  **
		"01100110", -- 8  **  **
		"01100110", -- 9  **  **
		"01100110", -- a  **  **
		"01111100", -- b  *****
		"01100000", -- c  **
		"01100000", -- d  **
		"11110000", -- e ****
		"00000000", -- f
		-- code x71
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01110110", -- 5  *** **
		"11001100", -- 6 **  **
		"11001100", -- 7 **  **
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01111100", -- b  *****
		"00001100", -- c     **
		"00001100", -- d     **
		"00011110", -- e    ****
		"00000000", -- f
		-- code x72
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11011100", -- 5 ** ***
		"01110110", -- 6  *** **
		"01100110", -- 7  **  **
		"01100000", -- 8  **
		"01100000", -- 9  **
		"01100000", -- a  **
		"11110000", -- b ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x73
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"01111100", -- 5  *****
		"11000110", -- 6 **   **
		"01100000", -- 7  **
		"00111000", -- 8   ***
		"00001100", -- 9     **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x74
		"00000000", -- 0
		"00000000", -- 1
		"00010000", -- 2    *
		"00110000", -- 3   **
		"00110000", -- 4   **
		"11111100", -- 5 ******
		"00110000", -- 6   **
		"00110000", -- 7   **
		"00110000", -- 8   **
		"00110000", -- 9   **
		"00110110", -- a   ** **
		"00011100", -- b    ***
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x75
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11001100", -- 5 **  **
		"11001100", -- 6 **  **
		"11001100", -- 7 **  **
		"11001100", -- 8 **  **
		"11001100", -- 9 **  **
		"11001100", -- a **  **
		"01110110", -- b  *** **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x76
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11000011", -- 5 **    **
		"11000011", -- 6 **    **
		"11000011", -- 7 **    **
		"11000011", -- 8 **    **
		"01100110", -- 9  **  **
		"00111100", -- a   ****
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x77
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11000011", -- 5 **    **
		"11000011", -- 6 **    **
		"11000011", -- 7 **    **
		"11011011", -- 8 ** ** **
		"11011011", -- 9 ** ** **
		"11111111", -- a ********
		"01100110", -- b  **  **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x78
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11000011", -- 5 **    **
		"01100110", -- 6  **  **
		"00111100", -- 7   ****
		"00011000", -- 8    **
		"00111100", -- 9   ****
		"01100110", -- a  **  **
		"11000011", -- b **    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x79
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111110", -- b  ******
		"00000110", -- c      **
		"00001100", -- d     **
		"11111000", -- e *****
		"00000000", -- f
		-- code x7a
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00000000", -- 4
		"11111110", -- 5 *******
		"11001100", -- 6 **  **
		"00011000", -- 7    **
		"00110000", -- 8   **
		"01100000", -- 9  **
		"11000110", -- a **   **
		"11111110", -- b *******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x7b
		"00000000", -- 0
		"00000000", -- 1
		"00001110", -- 2     ***
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"01110000", -- 6  ***
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00001110", -- b     ***
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x7c
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2    **
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00000000", -- 6
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"00011000", -- b    **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x7d
		"00000000", -- 0
		"00000000", -- 1
		"01110000", -- 2  ***
		"00011000", -- 3    **
		"00011000", -- 4    **
		"00011000", -- 5    **
		"00001110", -- 6     ***
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"01110000", -- b  ***
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x7e
		"00000000", -- 0
		"00000000", -- 1
		"01110110", -- 2  *** **
		"11011100", -- 3 ** ***
		"00000000", -- 4
		"00000000", -- 5
		"00000000", -- 6
		"00000000", -- 7
		"00000000", -- 8
		"00000000", -- 9
		"00000000", -- a
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000", -- f
		-- code x7f
		"00000000", -- 0
		"00000000", -- 1
		"00000000", -- 2
		"00000000", -- 3
		"00010000", -- 4    *
		"00111000", -- 5   ***
		"01101100", -- 6  ** **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11111110", -- a *******
		"00000000", -- b
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000"  -- f
	);
begin
	process(addr)
	begin
	data <= ROM(to_integer(unsigned(addr)));	
	end process;
	dataOut <= data;
end Behavioral;